`default_nettype none
module tt_um_noritsuna_8bitcounter (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

reg [7:0] count;
assign uo_out = count[7:0];
assign uio_out = count[7:0];
assign uio_oe = ena == 1'b1 && count < 8'b11111111;
always @(posedge clk) begin
        if (rst_n == 1'b0) begin
                count <= 'b0;
        end else if (ena == 1'b1) begin
                count <= count + 1'b1;
        end
end
endmodule
